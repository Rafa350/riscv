`ifndef __RV_SVH
`define __RV_SVH


// Model i extensions del procesador.
//
`define RV_BASE_RV32I
`define RV_EXTENSION_C
`define RV_EXTENSION_M

// Adresses dels vectors
//
`define RV_VECTOR_RESET  32'd0
`define RV_VECTOR_NMI    32'd4


`endif
