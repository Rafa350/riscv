module HazardDetector(
    output logic [1:0] o_DataASelect,
    output logic [1:0] o_DataBSelect);


endmodule
