module FPU
(
    );

endmodule
