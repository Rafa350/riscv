module FPU
    import CoreDefs::*;
(
    );

endmodule
