// -----------------------------------------------------------------------
//
//       Memoria de lectura/escriptura.
//
//       Lectura asincrona i escriptura sincrona.
//       Un canal per lectura, i un altre per escriptura.
//       Escriptura i lectura simultanies.
//       Es direcciona en bytes pero retorna word de DATA_WIDTH bits
//
//       Parametres:
//           DATA_WIDTH : Amplada del canal de dades
//           ADDR_WIDTH : Amplada del canal d'adresses
//
//       Entrades:
//           i_clock    : Rellrotge
//           i_addr     : Adressa per escriptura i/o lectura
//           i_wre      : Habilita l'escriptura
//           i_data     : Dades per escriure
//
//       Sortides:
//           o_data     : Dades lleigides
//
// -----------------------------------------------------------------------

module RwMemory
#(
    parameter DATA_WIDTH = 32, // Amplade de dades
    parameter ADDR_WIDTH = 32) // Amplada d'adresses
(
    input  logic                  i_clock, // Clock

    input  logic [ADDR_WIDTH-1:0] i_addr,  // Adressa
    input  logic                  i_wr,    // Habilita l'escriptura
    input  logic [DATA_WIDTH-1:0] i_data,  // Dades per escriure
    output logic [DATA_WIDTH-1:0] o_data); // Dades lleigides

    localparam SIZE = (2**ADDR_WIDTH)>>2;

    logic [DATA_WIDTH-1:0] data [0:SIZE-1];

    always_ff @(posedge i_clock)
        if (i_wr)
            data[i_addr[ADDR_WIDTH-1:2]] <= i_data;

    assign o_data = data[i_addr];

endmodule
