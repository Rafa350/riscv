`define RV_BASE_RV32I
`define RV_EXTENSION_C
`define RV_EXTENSION_M
