module FPU
    import ProcessorDefs::*, CoreDefs::*;
(
    );

endmodule
