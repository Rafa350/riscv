module MultDiv;


endmodule
