module stageE

endmodule
