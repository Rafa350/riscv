module Divider
    import Types::*;
(
    input Data i_operandA,
    input Data i_operandB);    


endmodule
