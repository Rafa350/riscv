module FPU
    import Types::*;
(
    );

endmodule
