module stageW(
);

endmodule
