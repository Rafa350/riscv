`define ALU_OP_A        4'h0
`define ALU_OP_B        4'h1
`define ALU_OP_AaddB    4'h2
`define ALU_OP_AandB    4'h3
`define ALU_OP_AorB     4'h4
`define ALU_OP_AxorB    4'h5
`define ALU_OP_notA     4'h6
`define ALU_OP_AeqB     4'h7
`define ALU_OP_AgtB     4'h8
`define ALU_OP_BshlA    4'h9
`define ALU_OP_BshrA    4'hA
`define ALU_OP_Ainc     4'hB
`define ALU_OP_Adec     4'hC

