module stageWB(
);

endmodule
