module StageWB();


endmodule
