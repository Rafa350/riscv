module pgm
#(
    parameter ADDR_WIDTH = 16,
    parameter INST_WIDTH = 16)
(   
    input  logic [ADDR_WIDTH-1:0] i_addr,
    output logic [INST_WIDTH-1:0]  o_inst);



endmodule