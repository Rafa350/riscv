module HazardDetector(

    output logic o_IFID_Stall,
    output logic o_IDEX_Flush,
    output logic o_EXMEM_Flush,
    output logic o_MEMWB_Flush);


endmodule
