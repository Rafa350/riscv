module stateM(
);


endmodule
